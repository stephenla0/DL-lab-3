module sevensegcall(
    a
);