module state_sel(
    a
);