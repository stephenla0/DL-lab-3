module top(
    a
);

