module sevenseg(
    a
);