module state_exe(
    a
);