module state_exe(
    output[2:0] state_select,
);